`include "ALUsync.v"
`include "clock.v"
module microprocessor(
  input wire [1023:0][7:0] memory, // Changed to wire to align with module instantiation
  input wire enable,              // Changed to wire
  output wire [7:0] result,
  output wire running
);

  integer file, code, t;

  reg [7:0] ar1, ar2;          // ALU's first and second register
  reg [7:0] arr;               // ALU's result register
  reg [5:0] operation_alu;     // ALU operation register
  reg [7:0] reader;            // Register to read bytecode
  reg enable_clk;              // Clock enable signal
  reg clk;                     // Clock signal
  wire fusion_enable = enable & enable_clk; // Combined enable signal
  wire alu_done;               // Signal indicating ALU operation completion
  integer line;                // Current line in the memory

  // ALU instance
  alu ALU (
    .clk(clk),                 // Connect clock
    .reset(enable_clk),        // Use enable_clk as reset
    .alu_start(enable),        // Connect enable as ALU start signal
    .a(ar1),                   // Operand A
    .b(ar2),                   // Operand B
    .op(operation_alu),        // ALU operation
    .result(arr),              // ALU result
    .alu_done(alu_done)        // ALU done signal
  );

  // Clock generator instance
  clock_gen CLOCK_GEN(
    .enable(fusion_enable),    // Enable clock generation when both enables are active
    .clk(clk)                  // Output clock signal
  );

  // Outputs
  assign running = enable_clk;
  assign result = arr;

  // Initialization
  initial begin
    enable_clk = 1;
    line = 0;
  end

  // Main operation logic 
  always @(posedge clk) begin
    if (alu_done)begin
    if (line == -1) begin
      enable_clk <= 0;         // Disable further operations
      $finish;                 // End simulation
    end else begin
      reader = memory[line];   // Read instruction
      $display("%b %b %b",result, ar1,ar2);
      case (reader)
        8'b00000010: begin     // Two-operand instruction
          line = line + 1;
          operation_alu = memory[line];
          line = line + 1;
          ar1 = memory[line];
          line = line + 1;
          ar2 = memory[line];
        end
        8'b00000001: begin     // Single-operand instruction
          line = line + 1;
          operation_alu = memory[line];
          line = line + 1;
          ar1 = memory[line];
        end
        8'b11111111: begin     // Termination instruction
          line = -2;           // Mark end of execution
        end
      endcase
      line = line + 1;         // Advance to next instruction
    end
    end
  end
endmodule
